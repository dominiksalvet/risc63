----------------------------------------------------------------------------------------------------
-- Copyright 2020 Dominik Salvet
-- github.com/dominiksalvet/risc63
----------------------------------------------------------------------------------------------------
